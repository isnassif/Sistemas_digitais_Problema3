module copia_direta (
    input clk,
    input reset,
    output reg [18:0] rom_addr,
    input [7:0] rom_data,
    output reg [18:0] ram_wraddr,
    output reg [7:0] ram_data,
    output reg ram_wren,
    output reg done
);

    parameter TOTAL_PIXELS = 160*120; // pixels da ROM

    reg [18:0] counter;
    reg [7:0] rom_data_reg;

    always @(posedge clk or negedge reset) begin
        if (!reset) begin
            counter <= 0;
            rom_addr <= 0;
            ram_wraddr <= 0;
            ram_data <= 0;
            ram_wren <= 0;
            done <= 0;
            rom_data_reg <= 0;
        end else begin
            rom_data_reg <= rom_data; // pega dado com 1 ciclo de atraso

            if (counter < TOTAL_PIXELS) begin
                rom_addr   <= counter;
                ram_wraddr <= counter;
                ram_data   <= rom_data_reg;
                ram_wren   <= 1;
                counter    <= counter + 1;
            end else begin
                ram_wren <= 0;
                done <= 1;
            end
        end
    end
endmodule
